`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 24.03.2024 09:48:09
// Design Name: 
// Module Name: mux
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux(
    input a,
    input s0,s1,s2,s3,
    output reg [15:0] y
    );
    
  always@(*)
   begin
     case({s0,s1,s2,s3})
     4'b0000:y={000000000000000,a};
      4'b0001:y={00000000000000,a,0};
      4'b0010:y={0000000000000,a,00};
      4'b0011:y={000000000000,a,000};
      4'b0100:y={00000000000,a,0000};
      4'b0101:y={0000000000,a,00000};
      4'b0110:y={000000000,a,000000};
      4'b0111:y={00000000,a,0000000};
      4'b1000:y={0000000,a,00000000};
      4'b1001:y={000000,a,000000000};
      4'b1010:y={00000,a,0000000000};
      4'b1011:y={0000,a,00000000000};
      4'b1100:y={000,a,000000000000};
      4'b1101:y={00,a,0000000000000};
      4'b1110:y={0,a,00000000000000};
      4'b1111:y={a,000000000000000};
      
      endcase
      end
      
                
            
endmodule
